`ifndef BRAM_PKG_SVH
`define BRAM_PKG_SVH

package bram_pkg;

    parameter LOW_LATENCY = 0;
    parameter HIGH_PERFORMANCE = 1;
    parameter NC = 0;
    parameter RF = 1;
    parameter WF = 2;

endpackage

`endif
